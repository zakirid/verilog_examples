module fa(a,b,cin,sum,co);
input 